//add primary io to system instance


   //CLINT
   input rtc,

assign rtc = rtc_in;

assign rtc = 1'b0;
